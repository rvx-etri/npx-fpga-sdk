`ifndef __MUNOC_PROCESS_ID_H__
`define __MUNOC_PROCESS_ID_H__

`define PROCESS_ID_I_MNIM_I_MAIN_CORE_NO_NAME (0)

`endif